module adder8(
        input  [7:0]  a,       //data in a
        input  [7:0]  b,       //data in b
        input  [7:0]  cin,     //cin
        output [7:0] sum_out,  //sum output
        output c_out           //carry output
        );
endmodule

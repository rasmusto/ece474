module testbench

module fifo (
);
